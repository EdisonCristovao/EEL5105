library IEEE;
use IEEE.std_logic_1164.all;

entity TOPO is 
port(

	A, B, C, D:in std_logic 	
);
end TOPO;

architecture circuito of TOPO is 

-- componentes


begin

end circuito;
